`ifndef SP_DEFAULT
`define SP_DEFAULT

// File included by SandPiper-generated code for the default project configuration.
`include "/home/shivani/Documents/self_study/test/out/sandpiper.vh"


`endif  // SP_DEFAULT
